package ahb_apb_test_pkg;

	import uvm_pkg::*;


	`include "uvm_macros.svh"

	`include "ahb_trans.sv"
	`include "ahb_agent_config.sv"
	`include "apb_agent_config.sv"
	`include "ahb_apb_env_config.sv"

	`include "ahb_driver.sv"
	`include "ahb_monitor.sv"
	`include "ahb_sequencer.sv"
	`include "ahb_agent.sv"
	`include "ahb_sequence.sv"

	`include "apb_trans.sv"
	`include "apb_driver.sv"
	`include "apb_monitor.sv"
	`include "apb_sequencer.sv"
	`include "apb_agent.sv"
	`include "apb_sequence.sv"

	`include "ahb_apb_scoreboard.sv"
	`include "ahb_apb_env.sv"
	`include "ahb_apb_test.sv"

endpackage

